//Объявление модуля универсального счетчика
module ucounter
#(
	parameter p_start_value = 0,			//Параметр отвечающий за начальное значение счета (нижнюю границу)
	parameter p_finish_value = 255		//Параметр отвечающий за конечное значение счета (верхнюю границу)
)
(
	input		logic		i_clk,				//порт сигнала синхро частоты
	input		logic		i_reset,				//порт сброса
	
	input		logic		i_set,				//порт управляющего сигнала установки начального значения
	input		logic		[def::numofbits(p_finish_value)-1:0] 	i_initial,	//Порт с начальным значением
																								//numofbits - функция, определенная и импортируемая
																								//из пакета def
	
	input		logic		i_work_enable,		//Порт разрешения работы счетчика
	input		logic		i_up_down,			//Порт определяющий направление счета
	
	output	logic		o_impulse,			//Порт выходного импульса по достижении крайнего значения
	output	logic		[def::numofbits(p_finish_value)-1:0]	o_data	//Порт выходного значения

);
	
	//Процедурный блок определяющий триггерную логику (ff - означает flip-flop, то есть триггер)
	//Все переменные блока работают по фронту (posedge) сигнала синхрочастоты (т.е. меняют свои значения только в
	//данный промежуток модельного времени и одновременно),
	//а также имеют ассинхронный сброс (наличие второго сигнала) по спаду (negedge) сигнала сброса
	always_ff @(posedge i_clk, negedge i_reset)
		//Часть кода описывает значения переменных во время асинхронного сброса
		if (~i_reset) begin
			o_impulse	<= 0;
			o_data		<= p_start_value;
			end
		//Часть кода, описывающая значения переменных при подачи сигнала установки	
		else if (i_set == 1) begin
			o_impulse <= 0;
			o_data <= i_initial;
			end
		else begin
			//Часть кода описывает работу счетчика при разрешающем сигнале работы
			if (i_work_enable == 1) begin
				//Описание работы инкрементного счетчика
				if (i_up_down == 1) begin
					if (o_data == p_finish_value) begin		//При достижении верхнего граничного значения
						o_data <= p_start_value;				//счетчик сбрасывается в начальное значение
						o_impulse <= 1;							//и устанваливается выходной импульс
						end
					else begin 
						o_data <= o_data + 1;					//В противном случае продолжается счет,
						o_impulse <= 0;							//а импульс или сбрасывается (чтобы он держался не дольше
						end											//одного такта), или находится в неактивном состоянии
					end
				//Описание работы декрементного счетчика	
				else begin
					if (o_data == p_start_value) begin
						o_data <= p_finish_value;
						o_impulse <= 1;
						end
					else begin
						o_data <= o_data - 1;
						o_impulse <= 0;
						end
					end
				end
			//Часть кода описывает поведение счетчика при запрещении работы
			else begin
				o_impulse <= 0;			//Выходной импульс устанавливается в 0
				o_data <= o_data;			//Значение счетчика не меняется
				end
			end


endmodule

